
module circuito(Us, Ua, H, T, M, L,Vs, Bs, Al, Cheio, Medio, Baixo, Critico, Erro, Ve);

always @(*) begin
   
end

endmodule
